PK   e{nWeF�i�'  w�    cirkitFile.json�ݎ�H��oŨ�����M�l�`g��Ә�6R$�%�J5��F_���^�fPeW�%�⍶w?��ۖ����`0�df�/W����\mwm��vw��n�^R��z[���O�������o˟v���W/�'��o�z�VM���.yQ�\ҭ�<�&���˻� �<�+��4��z�����-�؂)I� �`J+f�Z0�3H-�ҋ�L�	Az���W�w﷛v�/��6�6I��N|VI�fibVi����+J�d�/�7^�T���y��]��ַ��|���v��?��wB_ʮ�I��L��\���ї��'�/3�m��SC.l�L؞��
���N�����g���K��D��?w�&"���+6)��Bj"R�r
��H!M�$7)�iWl"R�SgoB�8��<�~y�M<��YH�@��{�6����Ek &X��@l"Rȟb�吘"Hc,@cL�l������ǒͤM�&њ�'6a8�)����Kb�B�h����AoB��"#����$�D�$��cIl"R�Kb�B�(�����D���p��H!��b����e�B:P���_l"R���D���l��Hx1#ϻ^�w�&"�<�MD
y����+6)�yWlA�w�&"�<w�MD
y�����)6)�Sl"R�s��D���N��H!ϝb�B�;�&"�<w�M�2��N��H!ϝb�B�;G&��<��QO�9ǐ�#,a�LIX��wP:�ҙ�b}g�����Δ�;�����tQC`}籾���.�!��X�A�K7�����)�Ax~tm0s�gب͆t���DI�k���\�c=�c�JGX:SX�X�A�KǓ_�s����������V6hi�67V7X>��Ti���
�G`>���X�`�������+,��xb=�`���#0/	 �گ'0��x1�`��#0����F�{�K*��{yt��c�`�b���G`��jY�Y�Y��_����W;�w;�;`�c��ǂ����|��	�?�����o�J�>�4}�����p� ��'OX>�/����s��.��_��]`�e���G`>^������|��<9,��|��5�`������|�+9!�����Y��{yt���BύCO�Cώ�'O,��|��%�`������|���?�������i��~u��#0/0�,_�|���`������|���?�/X>�qI�����G`>.� ������|\��?������P���^��^����˛��]��ōK����A\�.~$�ݔ��B�4:qiBW�U��,�����`Ճ�#0���z�|��:X����������V=X>�q#�����G`>.��X�`��ǥ����,���������`���%�ߺ`��ǅ����,���D�`���#0w��?�|��tX��`���#0���?�|��R�`�����.�-�փ\�W���aƅ���.���;1S���.�^ɠK'@�|]x��V��{�+Rɵ�6}\z��v"+�|�D�/�G{#.=_x��#\z�0�G{ .=Xbxi6��h�����ݖ�/�?+�W:H�Ѧi�7$�%oD�����/�m����{�:_8��ę&$>J��|�]��y�EE<��N���;����6wm�j�tYۮZuI�E�{O)���ՙk�u����:}��몰M�x��&�Ɋ$o�4�i�*ڦɫڜ��u�4��ӧ���eu�UҵM��̹$/r����M�W����>��@�M�le��>���E�g�MC�8����ӧ��4�\(SD��!���&m[�(\U�s7������/��r����^�"y|D��ߙ�����/O� C�Eb�@�����N~"�!úC2��h��
��2���w�ɉR�!:�_WC��(/~���e�V�Qq�c.��� �d��C���ڸ���K�(K�� 1�r7��7ʒ��e@L K��1�,�~����K�(K��1�'���񏖲�B&X?XB��,�����Q�L?	b��q�����<�`�����L�<nA�z����`y���8ʒ��qAr�w�<��ĕu`L�7��[��T]'d��q�%.�c���,��,q��?�`ye��L��`y�����RZ�6]	�`ye�K��`�q��(K������Q�x&�	��=,��,�"_,�{XGY�Ũ(&�%^�	c��� ��(K������Q�x��	��,��,��.,�XGY�H0&XOaye����`y<���)K�W�O����XVI��TXM9\W�
��+���r��
n�WVRa5��*Я���u��_�U"0�`%��R��z�����(#��\�U�_Ǭ`�@��L��>��ߵ-��+�`Ex`Xn����j�a]
�U�_5XI����ťBK:�<�YǷJ�KIv��.�^���ThI�����VG}�В-ϙ��S�%Z����[�BK:���AǷ:JL��thy-��o5�В-�)��"S�%Z^��۱�A�"���)Z���.�:�L��thy��ʠ���e'h�f��Uz!��FL镘�.�:����2Zҡ�5p:���e*��C�k�t�.;A�6����.�:�L��thym��ouޒ���)Z�tt���e*��C�k]u|��L��thyͮ��$]�BK:���XǷ:�L��thy��o�J�,S��S�'(MVT���4]QG�9]�tt�
-����|���2Zҡ�:���e*��C˵t|��L��th�惎out�
-��r�
���2Zҡ�*��:�L��th����out�
-��rM��/S�%Z���[]�BK:�\�FǷJ+ɔ�����^o��e^G���E�E�VG�7������)Z�tt���e*��C�5�t|���ThI��kQ��VG��В-��R�m��e*��C˵�t|���ThI��k���VG��В-�j��.S�%Z�9��[]�BK:�\;OǷJU>��|�負�˂��2Zҡ�Z�:���e*��C�5u|���ThI��kK��VG��В-��T�m���ThI��k}��VG��В-�,��.S��y�7���t���DmڅV&��.��bş~����D��V���Z��G���D�V5�G��-�:P�b�����xC��f0�;���R3����t�LOm���D��Y�S;q.5�I�S�T.5��b;���R3�(>�8��i�L��p��ҧ.&��v|4c�/�mm�L%yp>��$Wdm^wQ�^��e�r�e�����6_�uH�,�}�j�%yM�=����V��2��E�̲r�/uU�&�M���o�"��"Ml����i�6��h���W4���+�C���VI�6E�3璼�mRS7uk\��m4���+�m���&q�2��j��]�be�MC�8.�̲r���4�\(SDS��!�b�H�6FLQ���3Zz���,��f�����W����/�f�o��|��~��n��-�Ud�p�"���!2}^���^yB�@�L�b!D C�W�"�!ӫkȐ�:�d���B2d#���ڸ���K�(K�0P�a��n�%o�%s��0��7�8ʒ9.a�`9�`Ie���0L�<naye��0L��7�����Q��a������Q��aD�����Q��a������Q��a#�ay���8��_�1�FRpC)�<�`ye�����`y���8��e�1���q�%�c��q��(K\w�����Q����	7&���q��(K������Q�x�3�	��=,��,�z[ثX�<����;aL�<`ye��po7q�7ay<��8����1��x��q�%^gc�����Q�x]�	��SX���|��h��a)	�*���
�)G��V�~�`%VS��>�����J*��գ@[�U��TX��R�������A*~���x@��TXcEů�h��
�)G�'�V�~�`%VS�jO�����J*��՝@[�U��TXyN��0�Q\*��C�s�u|����d���"�E:�K��thy���ouԗ
-���y��(0Zҡ��:��Qa*��C�kt|���ThI���b��VG��В-�)��"S�%Z^��[U�BK:���G�ł�.S�%Z^���[]�BK:���JǷJoĔ^���2��ˬ�.S�%Z^��[]�BK:���OǷ:�L��thyM��out�
-����J���2Zҡ�5�:���e*��C�k]u|���ThI�����LL��e*��C�k�u|���ThI���P��VG��В-����lE��:����2���ThI������VG��В-���.S�%Z����[]�BK:�\�AǷ:�L��th�v��out�
-��r�z]�BK:�\KDǷ:�L��th�&��out�
-��rm���2Zҡ�5:�UZI���LG�y]�ut�
-��r� ���2Zҡ��G:���e*��C�5�t|���ThI��kQ��VG��В-��R�m��e*��C˵�t|���ThI��k���VG��В-�j��.S�%Z�9��[]�BK:�\;OǷJU>��|�負�˂�.S�%Z�e��[]�BK:�\�QǷ:�L��th����out�
-��r�Lߦ:�L��th�֧�out�
-��r�R���2Z�G�p/��J��LԦ]he���B+u�Z������D��V&�[/�2Q�z���
��L�|^u���D�Ԧ�K�`�wjkեf0<���R3���&t�LOmƹ�(c�xj�ʥf0Q<��R3�(��qq�LO�k��������X�g[�8ӄ�CI�Ob?�Y��]��afY��\��fY�x?��Wm�.�b�ZuI�ES�{O)����e�̲r�/��\�K]�I}�Am⛬H�H����m�����+�e��Ͳr���eu�UҵM��̹$/r����M�W�nFͱr�|���I��L��'u���FYgӐ5΄�,��\d�,+��є�|H��+���S��쌖�e�)˯��?����v�+���W/���>�w�]���Z�M�ޔ�]��^�z������SԵ|s-�y+��%tB���W�Kq�g��E�����Wg �ABg�Qr�p�Uˤ�1�����7�Q`>c�+�������d��C��"D��3F��ya��a�=M���%��R���u�엔���.�U#����곫7o>��w���cǼ�4���"h<�������C��=*���P�;�*a�������p�}^������Q#�@�G\Cb|%��(1ꖂ���� d2C��!rь��3�3>2��>r%}��3jRW����b�a��"�z�?x��l˻}�o�^~���������_7W/�$~�Y�'6qxE*��8�LR�M�~څ�Bl���Q�b���j����',�2�l�NY]��'�$#c�䍛�C,_��	��&�a��4!"�2"123R�܆9̔�r �3ҳ܆9�Ֆr�m��do)�؆9��r R+r�܆9�W�r�ǡh���K{zf�%i1���R,c�ơ�a~��|- ��m��
) �Z@�'��N����D�� �َ���
� �Zn��dH9 =_H�r�*D���:@��m�X�Q
7��7H�r�1��/v�\,�� 8 �bȶr\H�ȶ�m��#L�.�$_��m� �|= ��mp�l  �z@z���w� @z���*��5~����Un�k��9�6��*��O ��mp�N  �@>��ຐ @>�|*����| �Tn���8 �4�S���� ���O�6�������;�#0��L9��������|�վ�ك��G`>S����A���#0_�`������G`�ؿ �oT8\x�X>󍦥���&2q�g��QYp���`���.�Kc\��*���A��G`>S��}��A���#0O�Dw���LHhB���!\��E
Z�Z�Z��		M�p�>Dk0!�	y�0ڇh�&$4!O|F��Y���&�I�h��
��Є<��Cl�Є�&���h�
��Є�:0>�����h%?����t-[,Z��		M8.gs~i��>ƥh&�� 谄�m��nA��V1�b���&�U8h�U��Є�Bh���c\�5`B^��K�����$Ƈ��Q�NB�	`��Ǣ5��Є�D�C��0!�	yyz�	ZԀ		M�K�>D�0!�	��,c|8��\>�hQ3�z >�>�>�-jZ�8�����ޢ}�V1`BB�a��*LHhB^��!����Є�^�C�l��ך�}��-`BB�:y�=Z��		Mȋ��>D�0!�	� ڇ�/`BBr1��:LHhB.��!|�|�Z�K쏖�r�h�2ĸ-[����H�� L'��@��V1`BBrY��*LHhB.��!Zŀ		M��h�>h&$4!��A��b���&�2@h�U��Є\��C�����/�}�V1`BBr�(�����Ѳ%�eK@�m��Kv�}��)`BBr�1��:LHhB.���!Z��		M�e��>L�:LHhB.Q��!Z��		M����>D�0!]"\�������G%�n�)<T�u�޷���UX]�������FN�?*L����ByI���U�tb��^����^j@��Mٖ�F�x��F�o�f1i`��[j@�H��n-5 ��S]{��<����K�I�Ԟȧ���)���I��󅳭M�iB⃡$�'�+㊬��.*�3 �Η����f��gn�ܵ���C�eY��U�.ɳh�x�)�ַ�:w���?s���?s�uU�&�M�jj�dE��E��4]m��U}bo���u��<tYl�tmS$>s.ɋ�&�1uS���;��9���m���&q�2��j��]���Φ!k�	�~��g~��4�\(SD#��!����m���pUe϶߬�������y놷���x��9i���+�DqǛ{��c��ȕ���8�����g�E�;�}>&>��h�É�'>���g��6�a��gX>���ϰ|��3�S�>�r����}�'Ɠ���9q�xR<aN`�0'�NȺ<��5IWPl��1Q�F'z
Y�gl��ޚ�5�&iEx����h�U�q!+x3">��1���_�,�f�mQ%>6A�C�G�Ñ!>���k�US��&�c�&��5�4K��Ґ;ʫ$[�xaE���Dׅ�JkcW>�.���֛v�Q]�	��Owҳv�)�1I�D���K�ƄVHh3�p���I	�l/�Ƅ^J�
�8�@�y��=c�THH��pX�jL��M)��JaЦ��^�h�l*%o����,��R�/9���� ?H�3�%�c:+��ꖌߎC=;�[.�E�{fcIi^2���O:T���}y[��-���cu��v��n�=|E���Wv��{�ʍ��_��W��0�*}�*�?|���*�*F_��K��5ӧk_4}�h:q���w������mR�ޖO�a�����n��2+4�"�叻������>�]y�v{�q1

i��6�t���\]y�<E%�5Dm�]u{ז.���r����k���&�����Ga%SZ�j2_TE_r�#fn�.�$s�I�(Zf��}�o���?T�*Z������}�ۯ�^4�{�������n�[o8)m�w�o�������=���}r��o��*��������o�ݫ��0~y�����[׷��v�ܯwm�b����]�����~���<=�	ɮ�_o� ����z��*���Ik��:w�M��d�?Ɠ�Lo��c��`�̛�x�����m��y���zs��6��9�F&����ul���rՇ�j�[ݶ��*!{�6xV\� ��\��7���M|���Sg�SgdSg�Tv�v���Ӈ;����>*�s�*��J�����uZ�"Р!?~�҉/�����yt��o�}��{�4<~�>~ڷ��d�ǿ�'��[��q;<|1����#_?|>�.�������e߬�mww�;�n��Ƈ�4�����mM������4�|N{�s���J~��!�s�IO�^|��Ze�	m�غ��vU�IJչo
W�ì7k@sN�s~W�Ǐ��ޱ��<}ͳg����2���D%���.����鉨�(���WI��Eb#v���J���=�6�y�Q9k�|ֳ؍��~E�.��q��ជ��ԣ�_��·��܏���]��x��;���ÍӅ��S�w�B�xj���.f;j��Ub��j�4�����j�0�f�g�n�x2���b���a>���h.���x0�*����[�ћ�=�˧Fr�c����������_�v�&6i���j�S���\Q�RQ��c׼(������v7��������G"�'n���,w�k���#sC������n���?�?��:��[�����v�����7զ�;�7<��2A���Q�����!f��M]��"��&�E��qNO�̮���Һ�*~��fIU��i���*_�j�|�@��|�I56�Q���h��]p��z�����"�\�I2�J=�u[p����ɲ�l���e�P���{F�g�PBz�ǁ�K�kF_��l���/��점(��"�{jn\�F�����z������c/���*iҼMr_7m��A?��(lfM�xV؜��(��Q�={��� �~�Nۙf�x�c�7�v��n_|X�7�7�͋~��Ŷ{���#�(�>�Yy�>���O>y�e�_q6P����]�������տ��o����I�����~�m�7ͷ���Ӑ~����u��/�����W��+?�#���3t�<�1�f��	�<�N���_��ٞ����GFs�ڤ�'h�n��M�{����9�A�ț�&3!�!\�[���Y;���u�qO�y�=%o��E�PL���]�RWU>�
k��=?k��{�7�Q|����n�v�z���}���7/b��o_�ίw�oyw�q7��Igrk�-�g�4����q?�97�i�_���8���w��;�7}NZw��r��¦.����q�Y�}�ۤ�{q���/�^�Cu{[ݽ��{���ޑ_�H�I��16��e�o�4��"-(�2��q���/�~�*!�ވ���謽q�w.�r.�?�k~��r�
r6�J�8k}��V�k��m��+��C�;�꧞��J|Z�d�rn��f�6~�Χ�޶���37ia��?��Ǒu^�U�޶�7�����k���u�~����~����1WĀz}�����6U׽��~�C��7��M��h�Lo��4'�-^J���U�r�/������|��}���@���uLY��mo�ׯ__��������Y��?}���̞��)==�&��_��?�x�QdNv<�h�a����7����5�� �����xtL�31%^�c�R�a��\jg���A�	���mm��J3��?o�S��?�9�?8jn |�]�=8 6 ���(@P��K��
��R;�`Z�� )�SQ(�wZ�OQ<�y�q�n^�s�dw�Y���U�d�f���
)d���+f�s�<+���,����`1�^����)��!�慀�r���X���4����y��{Vs�AG"����a��a��ּ�}����ܨ���&��N'�Ӡ]���18l���
����G��������i)}HK��1��O玣���1�Q��B�gq!�й�,��*���0��ɨ��n.>��lC`�<7��"%z�rq����&n��y��f�R��=�>lf��̓GZ�F3�����0�������*=ж��FN��
l�S��_��D�H�~:ʆ�YZB	:颼�,Vd���ڝ�l�d��f����:�dMУ�ؿ��7��U��x�.t�O������s����M�ܦ+p�xd�dz������p�Θxy38jJ�Yj��
�������S�ow��7ډ�s��c��m�js_�~�}��}���u_�����PK   e{nWeF�i�'  w�            ��    cirkitFile.jsonPK      =   �'    